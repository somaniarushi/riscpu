`define RF_PATH   cpu.rf
`define DMEM_PATH cpu.dmem
`define IMEM_PATH cpu.imem
`define BIOS_PATH cpu.bios_mem
`define CSR_PATH  cpu.tohost_csr
