module alu (
    input [31:0] rs1,
    input [31:0] rs2,
    input [31:0] alu_sel,
    output reg [31:0] alu
);
endmodule