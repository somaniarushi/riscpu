module control_logic (
    input [31:0] inst_fd,
    input [31:0] inst_x,
    input [31:0] inst_mw,
    input brlt,
    input breq,
    // TODO: branch comparator input
    output reg [1:0] pc_sel,
    output reg is_j_or_b,
    output reg wb2d_a,
    output reg wb2d_b,
    output reg brun,
    output reg asel,
    output reg bsel,
    output reg alu_sel
);

    // Setting PCSel
    /*
        1. If the instruction in inst-FD is a JAL instruction, it's time to jump -> PC + imm, PC Sel = 0
        2. If the branch of inst-X is taken or inst-X is JALR, then jump to ALU value -> ALU, PC Sel = 1
        3. If none of the above 2 are true, go to PC + 4, PC Sel = 2
    */
    wire fd_is_jal, x_is_jalr, x_branch_taken;
    assign fd_is_jal = inst_fd[6:0] == 7'h6F;
    assign x_is_jalr = inst_x[6:0] == 7'h67 && inst_x[14:12] == 3'h0;
    assign x_branch_taken = 0; // FIXME: DO BRANCHING

    always @(*) begin
        if (x_is_jalr || x_branch_taken) begin
            pc_sel = 1;
        end else if (fd_is_jal) begin
            pc_sel = 0;
        end else begin
            pc_sel = 2;
        end
    end

    // Setting isJorB
    /*
        1. If inst-X is a JALR instruction, set to true.
        2. If inst-X is a branch instruction, set to true.
        TODO: Anything missing here?
    */
    wire x_is_branch;
    assign x_is_branch = inst_x[6:0] == 7'h63;
    always @(*) begin
        if (x_is_jalr || x_is_branch) begin
            is_j_or_b = 1;
        end else begin
            is_j_or_b = 0;
        end
    end

    // Setting wb2d-a
    /* Conflict between rs1 when rd of inst-MW = rs1 of inst-FD. */
    wire rd_instmw, rs1_instfd;
    assign rd_instmw = inst_mw[11:7];
    assign rs1_instfd = inst_fd[19:15];
    always @(*) begin
        if (rd_instmw == rs1_instfd) begin // a conflict exists, forwarding required
            wb2d_a = 1;
        end else begin
            wb2d_a = 0;
        end
    end

    // Setting wb2d-b
    /* Conflict between rs2 when rd of inst-MW  = rs2 of inst-FD. */
    wire rs2_instfd;
    assign rs2_instfd = inst_fd[24:20];
    always @(*) begin
        if (rd_instmw == rs2_instfd) begin
            wb2d_b = 1;
        end else begin
            wb2d_b = 0;
        end
    end

    // Setting brUN
    /* Branch unsigned = 1 if the inst type is B and func3[3:1] == "11" */
    wire x_is_unsigned = inst_x[14:12] == 3'b110 && inst_x[14:12] == 3'b111; // BLTU or BGEU
    always @(*) begin
        if (x_is_branch && x_is_unsigned) begin
            brun = 1;
        end else begin
            brun = 0;
        end
    end

    // Setting ASEL
    /*
        ASel = 0 when RS1 is used.
        ASel = 1 when PC is used. Instruction is AUIPC, or jump or branch
        ASel = 2 when WB forwarding is used. Conflict between rs1 and rd.
    */
    wire rs1_instx = inst_x[19:15];
    if (rd_instmw == rs1_instx) begin
        asel = 2;
    end else if (inst_x[6:0] == 7'h17 || inst_x[6:0] == 7'h6F || inst_x[6:0] == 7'h63) begin
        asel = 1;
    end else begin
        asel = 0;
    end

    // Setting BSEL
    /*
        BSel = 0 when RS1 is used.
        BSel = 1 when IMM is used. If the instruction is not an R-type, select IMM.
        BSel = 2 when WB forwarding is used. Conflict between rs2 and rd.
    */
    wire rs2_instx = inst_x[24:20];
    if (rd_instmw == rs1_instx) begin
        bsel = 2;
    end elif (inst_x[6:0] != 7'h33) begin
        bsel = 1;
    end else begin
        bsel = 0;
    end


    wire x_opc = inst_x[6:0];
    wire x_func3 = inst_x[14:12];
    wire x_func7 = inst_x[31:25];
    // Setting ALUSel
    /*
        ADD = 0, SUB = 1, SLL = 2, SLT = 3
        SLTU = 4, XOR = 5, SRL = 6, SRA = 7, OR = 8,
        AND = 9
    */
    // For R-Type
    if (x_opc == 7'h33) begin
        case (x_func3)
            3'b000: alu_sel = (x_func7 == 7'b0) ? 0 : 1;
            3'b001: alu_sel = 2;
            3'b010: alu_sel = 3;
            3'b011: alu_sel = 4;
            3'b100: alu_sel = 5;
            3'b101: alu_sel = (x_func3 == 7'b0) ? 6 : 7;
            3'b110: alu_sel = 8;
            3'b111: alu_sel = 9;
            default: alu_sel = 0;
        endcase
    end
    // For I-Type instructions
    else if (x_opc == 7'h03 || x_opc == 7'h13 || x_opc == 7'h67 || x_opc == 7'h73) begin
        case (x_func3)
            3'b000: alu_sel = 0;
            3'b001: alu_sel = 2;
            3'b010: alu_sel = 3;
            3'b011: alu_sel = 4;
            3'b100: alu_sel = 5;
            3'b101: alu_sel = (x_func3 == 7'b0) ? 6 : 7;
            3'b110: alu_sel = 8;
            3'b111: alu_sel = 9;
            default: alu_sel = 0;
        endcase
    end
    // For every other instruction -> default to add
    else begin
        alu_sel = 0;
    end

endmodule