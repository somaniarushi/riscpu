module immediate_generator (
    input [31:0] inst,
    output [31:0] imm
);
endmodule